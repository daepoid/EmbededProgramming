module bit_shift_blocking(A, B, C, D, E, clk);
  output A, B, C, D;
  input E, clk;

  reg A, B, C, D;

  always @(posedge clk) begin
    A = B;
    B = C;
    C = D;
    D = E;
  end
endmodule

